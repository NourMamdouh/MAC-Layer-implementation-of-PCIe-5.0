module phy_top #(
  serdes                       = 0,
  DATA_WIDTH                   = 256,
  BUFFER_DEPTH                 = 8,
  ADDR_WIDTH                   = 3,
  PACKET_LENGTH	               = 'd11,    
  SYMBOL_PTR_WIDTH             = 'd5,					
  SYMBOL_NUM_WIDTH	           = 'd4, 								
  SYMBOL_WIDTH		             = 'd8,           		  	
  MAX_LANES			               = (2**SYMBOL_PTR_WIDTH),
  FILTERED_Buff_DATA_In_WIDTH  = 30,
  FILTERED_Buff_DATA_Out_WIDTH = 31,
  FRAME_DEPTH                  = 4,
  SYNC_WIDTH                   = 2,
  BUFFER_WIDTH_ELSTC_BUFF      = 13,
  PTR_WIDTH                    =4,
  DEPTH_ELSTC_BUFF             =8,
  THRESHOLD_PTR_ELSTC_BUFF     =2,
  BITS_COUNT_WIDTH             =3
)(
  input                                   CLK,
  input  logic                            rx_clk, rx_rst,
  input  logic [0:DATA_WIDTH-1]           rx_data,
  input                                   RST_L,
  input                                   i_EN,
  input  logic                            GEN, 
  input  logic                            i_EN_BA,
  input	    							                i_Lanes,   			// 32 lanes or only one lane
  input                                   i_RD_EN,
  input [0:MAX_LANES-1]                   PIPE_d_K,
  // general outputs    
  input                                   i_EN_PF,
  input  [0:MAX_LANES-1]                  RXValid,
  input  [0:MAX_LANES-1]                  RX_Data_Valid,
  input  [0:MAX_LANES-1]                  RX_Start_Block,
  input  [0:SYNC_WIDTH-1]                 RX_SYNC_Header [0:31], 
  input  [1:0]                            i_GEN_Lanes,
  input                                   i_Os_Enable,
  input [0:(SYMBOL_WIDTH*MAX_LANES)-1]	  i_OS,
  input                                   i_WR_EN,
  input                                   i_SOP,i_End_Valid,i_Type,
  input [PACKET_LENGTH-1:0]               i_Length,
  input [SYMBOL_PTR_WIDTH-1:0]            i_Last_Byte,
  input [0:DATA_WIDTH-1]                  Data_IN,
  input                                   idle_cnt_enable,
  input [0:MAX_LANES-1]                   o_D_K,
  input                                   Soft_RST_blocks,
  input                                   type_IDL_TS,
  input                                   PIPE_CNT_rst,
  input                                   IDL_rst,
  input                                   rst_BA,
  output [0:MAX_LANES-1]                  back_pressures,
  output                                  ack_done,
  output                                  o_Full, // re consider the throttling of DATA LINK Layer
  output [0:(SYMBOL_WIDTH*MAX_LANES)-1]	  out_data, // GEN 3 
  output [0:MAX_LANES-1]                  valid_data, // GEN3
  output [0:MAX_LANES-1]                  TxStartBlock,
  output [0:1]                            TxSyncHeader [0:MAX_LANES-1],
  output    							                o_Idle_Indicator,  //raised one when sending idles (no more TLPs or DLLPs to send)
  output	    							              RX_Error,  				//to be raised when an error is detected
  output                                  o_Empty,
  output [0:DATA_WIDTH-1]                 Data_Out,
  output                                  o_SOP,o_End_Valid,o_Type,
  output [PACKET_LENGTH-1:0]              o_Length,
  output [SYMBOL_PTR_WIDTH-1:0]           o_Last_Byte,
  output [SYMBOL_NUM_WIDTH-1:0]           deskewed_RX_count [0:MAX_LANES-1],
  output                                  valid_deskew,
  output [0:DATA_WIDTH-1]                 Des_Data_Out,
  output [0:MAX_LANES-1]                  Block_Type,
  output                                  EIEOS_Flag,
  output                                  o_Sync_Sel
);

logic [0:MAX_LANES-1]                  BA_error;
logic                                  Deskew_error;
logic                                  PF_Error;

assign RX_Error = (Deskew_error | PF_Error | (|BA_error));

PHY_TX  #(
  .BUFFER_DEPTH(BUFFER_DEPTH),
  .ADDR_WIDTH(ADDR_WIDTH),
  .serdes(serdes),
  .SYNC_WIDTH(SYNC_WIDTH),
  .SYMBOL_NUM_WIDTH(SYMBOL_NUM_WIDTH),
  .SYMBOL_WIDTH(SYMBOL_WIDTH)
) u_PHY_TX (
  .CLK(CLK),
  .RST_L(RST_L),
  .i_EN(i_EN),
  .i_GEN_Lanes(i_GEN_Lanes),
  .i_Os_Enable(i_Os_Enable),
  .i_OS(i_OS),
  .i_WR_EN(i_WR_EN),
  .i_SOP(i_SOP),
  .i_End_Valid(i_End_Valid),
  .i_Type(i_Type),
  .i_Length(i_Length),
  .i_Last_Byte(i_Last_Byte),
  .Data_IN(Data_IN),
  .o_Full(o_Full), 
  .out_data(out_data), 
  .valid_data(valid_data), 
  .TxStartBlock(TxStartBlock),
  .TxSyncHeader(TxSyncHeader),
  .o_Sync_Sel(o_Sync_Sel),
  .back_pressures(back_pressures),
  .idle_cnt_enable(idle_cnt_enable),
  .ack_done(ack_done),
  .o_D_K(o_D_K),
  .Soft_RST_blocks(Soft_RST_blocks), 
  .IDL_rst(IDL_rst),  
  .o_Idle_Indicator(o_Idle_Indicator)  
);

PHY_RX #(
  .SYMBOL_WIDTH(SYMBOL_WIDTH),				          
  .PACKET_LENGTH(PACKET_LENGTH),				          
  .SYMBOL_NUM_WIDTH(SYMBOL_NUM_WIDTH),			        
  .SYMBOL_PTR_WIDTH(SYMBOL_PTR_WIDTH), 			       
  .MAX_LANES(MAX_LANES),					           
  .FILTERED_Buff_DATA_In_WIDTH(FILTERED_Buff_DATA_In_WIDTH), 	
  .FILTERED_Buff_DATA_Out_WIDTH(FILTERED_Buff_DATA_Out_WIDTH), 	
  .FRAME_DEPTH(FRAME_DEPTH),                   
  .DATA_WIDTH(DATA_WIDTH),                    
  .BUFFER_DEPTH(BUFFER_DEPTH),                  
  .ADDR_WIDTH(ADDR_WIDTH),                    
  .serdes(serdes),                        
  .SYNC_WIDTH(SYNC_WIDTH),                    
  .BUFFER_WIDTH(BUFFER_WIDTH_ELSTC_BUFF),                  
  .PTR_WIDTH(PTR_WIDTH),                     
  .DEPTH(DEPTH_ELSTC_BUFF),                         
  .THRESHOLD(THRESHOLD_PTR_ELSTC_BUFF),                     
  .BITS_COUNT_WIDTH(BITS_COUNT_WIDTH)              
) u_PHY_RX (
  .CLK(CLK),
  .RST_L(RST_L), 
  .rx_clk(rx_clk), 
  .rx_rst(rx_rst),
  .i_EN_BA(i_EN_BA),
  .rx_data(rx_data),
  .GEN(GEN), 
  .deskewed_RX_sync(Block_Type), 
  .EIEOS_Flag(EIEOS_Flag),  
  .Soft_RST_blocks(Soft_RST_blocks),  
  .type_IDL_TS(type_IDL_TS), 
  .PIPE_CNT_rst(PIPE_CNT_rst),
  .i_Lanes(i_Lanes),
  .i_RD_EN(i_RD_EN),
  .i_EN_PF(i_EN_PF),
  .enable_LDS(i_EN_BA),
  .PIPE_d_K(PIPE_d_K),
  .RX_Data_Valid(RX_Data_Valid),
  .RXValid(RXValid),
  .RX_Start_Block(RX_Start_Block),
  .RX_SYNC_Header(RX_SYNC_Header),
  .BA_error(BA_error),
  .Deskew_error(Deskew_error),
  .o_Empty(o_Empty),
  .Data_Out(Data_Out),
  .o_SOP(o_SOP),
  .o_End_Valid(o_End_Valid),
  .o_Type(o_Type),
  .o_Length(o_Length),
  .o_Last_Byte(o_Last_Byte),
  .PF_Error(PF_Error),
  .deskewed_RX_count(deskewed_RX_count),
  .Des_Data_Out(Des_Data_Out),
  .valid_deskew(valid_deskew),
  .rst_BA(rst_BA)
);


endmodule
